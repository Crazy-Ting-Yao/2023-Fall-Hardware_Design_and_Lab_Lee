`timescale 1ns/1ps
`include "Universal_Gate.v"




module Decode_And_Execute(rs, rt, sel, rd);
input [4-1:0] rs, rt;
input [3-1:0] sel;
output [4-1:0] rd;

endmodule
